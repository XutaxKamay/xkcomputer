library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.CentralProcessingUnit_Package.all;

entity CentralProcessingUnit is
    port
    (
        reset: in boolean;
        commit_read_memory: inout boolean;
        commit_write_memory: inout boolean;
        memory_size_read: out MEMORY_INTEGER_SIZE_TYPE;
        memory_size_write: out MEMORY_INTEGER_SIZE_TYPE;
        memory_address_read: out CPU_ADDRESS_TYPE;
        memory_address_write: out CPU_ADDRESS_TYPE;
        memory_data_read: in MEMORY_BIT_VECTOR;
        memory_data_write: out MEMORY_BIT_VECTOR
    );
end CentralProcessingUnit;

architecture CentralProcessingUnit_Implementation of CentralProcessingUnit is
    signal signal_reset_request: boolean;
    signal signal_unit_state: UNIT_STATE := UNIT_STATE_NOT_RUNNING;
    signal signal_registers: REGISTERS_RECORD;
    signal signal_has_asked_instruction: boolean := false;
    signal signal_memory_to_commmit: COMMIT_MEMORY_RECORD;
begin
    -- Handle control unit reset --
    process (reset)
    begin
        if reset then
            signal_reset_request <= true;
        else
            signal_reset_request <= false;
        end if;
    end process;

    ----------------------------------------------------------------------------
    -- Handle control unit states
    -- Feedback loop based on signal_unit_state FSM
    process (signal_reset_request, signal_unit_state)
    begin
        -- Reset has been raised --
        if signal_reset_request then
            -- Reset CPU --
            signal_registers <= (general => (others => (others => '0')),
                                 special => (overflow_flag => false, 
                                             condition_flag => false,
                                             program_counter => (others => '0'))); 
            -- In case we interrupted while being in commiting state --
            signal_memory_to_commmit.has_commit <= false;
            -- Do not wait for memory to set them to false --
            commit_read_memory <= false;
            commit_write_memory <= false;
            -- Will trigger again a new process execution --
            signal_unit_state <= UNIT_STATE_BEGIN;
        end if;

        case signal_unit_state is
            -- Should never happen --
            when UNIT_STATE_NOT_RUNNING =>
                signal_unit_state <= UNIT_STATE_BEGIN;

            -- This is an extra step, but maybe not needed, this in case we need extra logic --
            when UNIT_STATE_BEGIN =>
                signal_unit_state <= UNIT_STATE_FETCH_AND_DECODE_AND_EXECUTE;

            when UNIT_STATE_FETCH_AND_DECODE_AND_EXECUTE =>
                FetchAndDecodeAndExecuteInstruction(commit_read_memory,
                                                    commit_write_memory,
                                                    memory_size_read,
                                                    memory_size_write,
                                                    memory_address_read,
                                                    memory_address_write,
                                                    memory_data_read,
                                                    memory_data_write,
                                                    signal_registers,
                                                    signal_has_asked_instruction,
                                                    signal_unit_state,
                                                    signal_memory_to_commmit);

            when UNIT_STATE_COMMITING_MEMORY =>
                CheckCommitMemory(signal_memory_to_commmit,
                                  signal_registers.general,
                                  commit_read_memory,
                                  commit_write_memory,
                                  memory_data_read,
                                  memory_data_write,
                                  signal_unit_state);
        end case;
    end process;

end CentralProcessingUnit_Implementation;
    
