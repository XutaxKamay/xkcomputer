library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.CPU_Package.all;

entity CU is
end CU;

architecture CU_Implementation of CU is
begin
	process (all)
    begin

	end process;
end CU_Implementation;
