library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.CentralProcessingUnit_Package.all;

entity MemoryRead is
    port
    (
        address_in: in CPU_ADDRESS_TYPE;
        request_size: in CPU_ADDRESS_TYPE;
        value_out: out std_logic_vector((INSTRUCTION_SIZE - 1) downto 0);
        done_job: out std_logic
    );
end MemoryRead;